/*********************************************************************************************************************************
 * Name                 : typedefs.sv
 * Creation Date        : 21-03-2022
 * Last Modified        : 21-03-2022
 * Author               : Badam Mayur Krishna
 * Author's Email       : mayurkrishna.b@alpha-numero.tech
 * Description          : Typedefs for all assignment questions
 **********************************************************************************************************************************/

typedef bit[9:0] b10;
typedef bit[8:0] b9;
typedef bit[7:0] b8;
typedef bit[6:0] b7;
typedef bit[5:0] b6;
typedef bit[4:0] b5;
typedef bit[3:0] b4;
typedef bit[2:0] b3;


`include "async_fifo.sv"
`define WIDTH 8
`define DEPTH 16

module top
(reg [`WIDTH-1:0] din,
reg wr_en,
reg rd_en,
reg clear,




endmodule





module adder(
input a,b,ci;
)
begin

end

module testbench();
reg a;
wire b;
integer c;
logic d;
real e;
bit f;
byte g;
int h;
shortreal i;
time j;
initial begin
 $display("Default values: %b, %b, %b, %b, %b, %b, %b, %b, %b, %b",a,b,c,d,e,f,g,h,i,j);
end
endmodule

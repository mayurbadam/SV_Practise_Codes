module str;
string a="mayur k";

initial begin
$display("%0d",a.len);
end
endmodule

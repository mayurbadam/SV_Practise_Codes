module datatypes1;

input wire a, b;
output s, c;






endmodule

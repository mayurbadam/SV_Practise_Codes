/*********************************************************************************************************************************
 * Name                 : top.sv
 * Creation Date        : 21-03-2022
 * Last Modified        : 21-03-2022
 * Author               : Badam Mayur Krishna
 * Author's Email       : mayurkrishnamk@gmail.com
 * Description          : Top file for d-flipflop
**********************************************************************************************************************************/

module top;

endmodule

class environment;
endclass

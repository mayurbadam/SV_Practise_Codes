module uvm;
   import uvm_pkg::*;
   import hello_pkg::*;

   initial run_test("hello_test");
endmodule

class face;
int eyes =2;
string colour = "Grey";

endclass


class transaction;
DIN[N:0]
WR_EN
WR_CLK
RD_EN
RD_CLK
clear
FULL
endclass

/*********************************************************************************************************************************
 * Name                 : .sv
 * Creation Date        : --2022
 * Last Modified        : --2022
----------------------------------------------------------------------------------------------------------------------------------
 * Author               : Badam Mayur Krishna
 * Author's Email       : mayurkrishnamk@gmail.com
----------------------------------------------------------------------------------------------------------------------------------
* Description          : 
**********************************************************************************************************************************/

module dut (
            input  wire clk,
            input  wire req,
            input  wire reset,
            output reg  gnt
           );
  always @ (posedge clk)
  begin
    gnt <= req;
  end
endmodule 

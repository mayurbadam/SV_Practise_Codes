module streaming;
logic [31:0] a,b,c,d,e,f;
logic [95:0] A;

initial begin
	A=1;

	A = {	
end
endmodule
